XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����kF���`fa.���p4����q:�0�%RO;��h�;'bE������zv1��n�R�}At4r�-��ܯ��}y��TМx���(�&�S�˗��+�B9y٣dn<O��[��
�a�}���G�Ȫ��1>\*��7H;ڽ��B�K=�҄Q3�\��������
t��a�_=}�Б8Е�j�&۰��aaR��$���+pl$#�5=�ۃĢ=~�c�K�D���\���ɸ{
�������AN
�$Z�q���>���q'�Ql��[@�pI��Z��or�U���^��;�9���
�}mQ�Grx���k��n��x2/" ���>�Ӿ���US嘁v�G_AQ���ֳ�GjC,+OPs�#�

�4�#���t`�6��}�x�oޔ�f��
A�wk���Q��D��:���}�kB���^px����>��%���c]u�A�	�a� �h����O�o�!D�Rk�˒�O�p��Ĉ_�Ű;�Y�c�K�7=�g}�J�����z3�����oM��a+L��eiZl�|�H�;#&�Z�s2��� �o��[��T��0��7�[_�(��mFd���+��5����_D��|�z4Z�A���s7*�;8��ʏ���0M�� �Ɍ���4"���:l�̀41��NJ�ە�Ҙ]��yH�2�䠰��������P��H�����=�v��!��r�p��(_���:��NaLb<~eM��Oh]q�����E���Kޫ�k�XlxVHYEB     400     130�y��%U�����0�"h�R �+��\`~.�OJ�$�sF'V5)w����iL�[+���˹�:>z��s�gk�7sɲ�"��.�ڻ0��}��履
nTd�5��Eoi���	��_�{�i�8�\�]���X.��K�}�2����*���@����}��q�~l��U�$��-�z��
�!a���X��� �cq�Y3U�ݯ��j�`%h���~���9�z��� �>�\�4�����O�gY�[W�|SY:��^�J�@�,�
^�?��x��	���Uà�I�����F�~�w( �i�XlxVHYEB     400     180��}�=�OcN!�0��p��#7e)�aj�}VX9{���^�:��8��XT3�F������ߤU=�~C`Z����/��X�X3�68å��A� ���d:d�xh,u-K�E��d��+��~�_MJ�=&�P���n�_�K����<�C)A�����
������G'z�,�84ʸ�1���dfM7M�^D���4�U��`�.�e�Gx���4��qe�}��EqFj�M�QJ%��Cl8��YֶS��	�S��F�4�����.).��G?�+�k�'�ǒ�;��&|1(�G�P@*�C��ri����2����>�1�����w²�3UfS.���NC��я�M��i�s￈���Ւ�k�� \���<�-XlxVHYEB     400      e0��o���cq�����a٭��x7ˎ	�f����G��C��ٞB1z��P���:�����UM7��T�(F%����D������<z�U,I�NN��\\����п�YF��'MT�<0L?"���[#�"O4#��-��P�v�?l�,�yY�_�I���Ȭ�6�c��:�P�g�_���5�6{h2ȐJC�!���x��4������6�Zg���XlxVHYEB     400     130���1���
��W��iu��[Z�ـ#^Ol�=R�ok�Xo�o��P(�WwW����_?��sܩ]XNP�I�ߠ�ـ�FZ�S]+���D��{w��qh�l��
��<����ۆ��a�lE9�i������䐣�p۾�|D��B\$n;��7���䜆��>�d���9���J�^Ʃ����\K�
�|�YTu,~*�f��q�K6<�������6������q�x��N��KC�ff���m�e�6c���^�>��獀}���3�d#�3��l��BP������d��{��f��-�yXlxVHYEB     400     110i��9!.ʬ��2aX��ҌC}�iE{,�|���H�tF�=-��%=!��厣���)�2��R�э��~`%C������9��2�\ݐ����|G�G��ۨ�}��K,���>�K��7�[����'X "�Ys[`t�$�f��S�?y��An�{�e���Ҥ�CV�2ns�x]�b���ĀdG�K��-�'��$5�`):t!��d변�ñc��&9��G��i�ſ���t����I�(|�/!QJ��/����XlxVHYEB     400      f0��ƚ��9R}�n���	|�y*`ծ�+r��)��ƀ�x�������B�q��	-5Qds���9I��D�i'�x����
r;���ݧ=��Υc�Ι����� oM?>k�i�HC�b�;��zN�Am���s;����d�9���������j�?F
)T�m��6�����%?Qc���H�8)���1�L���ל'��-I���+J�����������nX&��i�"Te���hAXlxVHYEB     400     180� ����Yp�+�/�A����GL!B�����ɿS4����x��B���=}�mXEAt�[fVz�������z)'h)�>+�H-C��2�Pu�Hz�J�sX�hYW�s%��ӹ�[Pv��	n��"]���_��	�"�������fU�:xm�Ƥ[��W�� h����>�nS[X��4U�{O�}t
G;��,��U�%�#f/��!���|�Fn�W,W��P���b�7��ymt�/�\0��MS�Ŀ�1��Fv����JԞ@f�ՈS�nE�ˊ�@ߗ����~�������/�8�y�� �Ղ챲�q�Y{{Zm��}��9r�k\?�(&��+.>]M�-��=��t7��u{��L~G�&�QcS\�dpXlxVHYEB     400     110��^������ 0;�{��"�>�I�Y���L�F�M@y�B���6��e䛴�l�����/���3��}��h�&q�tCܼ6 (qEN�S�1y������D�zFð*7�ݦ�3��G��h^�o$H���N�N����'����teO�*6K���&�H�����޼<'~��+�����j�R��gx� �H�w���DL����o��ZZ(:
E��p<�3�aX����jV,�w�v�� �	_��^n~�O���w�ی2VXlxVHYEB     400     150�wl��6��E!��%h��ʙ���j?��yV^����t^wd�ihw	�}5:�[Qk�a-� ���?n� kt�Ab�����X[L��ޖ�v�6���AJD�d��e��Zل���Uf#X����5�S�@�Ԝ���k���p�&���RS#�Ĭ��A��%�̘�	�МI�"7 w$nu�
��8s����.œf�ȇ`����"��B�[���r۽}{v�Ѱp��*Z��1�0Zl�n�M`����ڵ��e�v��WfF�P�D��f���޶Lq&;~3����h���� �O"W�9n�K�^)����s��Y�~��%����E�XlxVHYEB     400     150�ssQ�&�Le`# ;V6��ӷD�'>�=����4� ��rXQ�%�~��S���Lu���O�͂�UB��xs�n���y�������GҶ�q�������{g{��H?0Y��{�Bu�"H�q�W��'�B�S�N�0`�V�7y����}q��nĪ�ڏ��.�Yx�(��T��ʏR����O�p�=�����GR�a���$d��?��"Рi���Z9�����@��:FB?i�V�M��Yl�*�C\+��P&E�ڢ
jߎ�kC�Ox����g=�>e�)��SBn0��LR5���>��f�m�{r(~�#fCcTz<iň���8�XlxVHYEB     400     110P�7Bw��:����{h$p�gE���'��yc���F��< ��ȁ8Q�s �=(�VN(�zc�r�����[N��t�A�����&���Kn� �_i}�̬�E��t��i�}I����u��A;X�*�������� j;<j���pPp���%+�uo�Rs�{��骬uGT���e�f,K&&c~fM鯎Ʈ�v�
�-𺇠��;��<�$��e���&1�]����QK��^�ȓt��r�5���8XJ|+�Z��bXlxVHYEB     400      a0���3djټ'��Zwy���%>��#؜g�Q�e��轉i�.qj�����-���\�;���~���(l_7��AɜW�ޭ��bم�Q��<Y��0n爷�Mm<�;��y�����X��_���,�{@����61�,#���J"�/��������XlxVHYEB     400     1d0��m�U,/�{Vg�m��x{�ת�T!���3ba����ك���Б�h�\����C���?2KSܫ�-s�S�{C<'څ�9Uo�M��DX)�;����sFe�h�Ȉ<�X�'":A+�r�d4"e,?�7㈑qZe��^k�m�����]�x�߶��V �r[��s�@m�*�.��x%�"�%��iM�<�Q�G�P~��#ͨNJ-��V\e�|��}u4f�_�19"��N`@�v��)�oDw�M��v�m�N�*���bT�/�[\�����&[uJY�5�_�XF����ݨ���g�e�~��T�Q�5��H5���P,M3@v 0T˛̳	���Κ�Y��U���&2B��eQ;�����\i���[dB4`���yq�`|ꁰrØ���;�+����1{bC�L��7�f1��A�"<m�_9/g�8;)�R@iTU���p���#�IE8XlxVHYEB     400      d0�r>�0������9YP1�����B;�!� )JuūY P�!*l��
4
����ʬܮ�?�1=JG��2ڈ�|C�?d-��ג%E�w�����h��J'aȮI����t���:�������O9�:icq�m
�G� {�D+���������z	.�Sk�p��ݽv\�l�Q#�_ZO�S*O�(�_��}:��fY8U�h٦��-bXlxVHYEB     400     130[�,���Cn:;�Q�Iߙv<��!�:������a���:g=Yh�KԾ������H�Q��Sk�G��XE����� v�D�O
p)��7����X>�'������O�U��C�H�mI�����'2��_�X�m����Je�� �	Q4�6�`J#�Qv��l�a?J�G�(o������k���S(P��ݰ�#Ҏ���y-n�f���5���:0Oکg�D�7B�!/�nֲnL�]8>=r���j��Ӿ�ں���X��wR�H����x�蒲�H��;u[�ja�銢P�I�B�0@B�BXlxVHYEB     400      b0��8�ž�N��eM���Ja�|Alغ˒�H���q�3�£�����#]�ϵ���W�;Wh�+u�[��V��fJ��3��	?{)�Z!5�_Y�l2"p�I�3*��(�
n�����U�81��`ΐ��UR*{z�8*V��k�dn���5?<���4�������:�X��8N,XlxVHYEB     400      f0���
ʁl��[ׂ�(ð���q�Ҙ�i>�,����N�բM�5:T��ł���&�Z�}�|"�t�mg���}L�|��� ���B9�Kb7�\=l۽h$r��>�TL��|^��}hV��	�l�U)-���,�F���22��X� �=�uN˯��!F�l��X��e��q}!�F�©J��b�$�Y�{��$�x�ӛC�%q���u�"v�诶ةiGϝ�w�:���I�XlxVHYEB     400      e08Z����ɱ�.)䝨J�|���/ʐQ�I�T����&�0�'~"_��̧�aQ�C��D,3��9+�O_�6C_�X���xY	+����$ �£��q��;�عoKg��������r�N��U�4	��n���:�~�_�l��ˋO���7{<Mj�_����nN�U�¹?6��'��� ct!&�����%ۯ����<�K�>�0�+x�XlxVHYEB     400     190���bA~i�V�%̺�P���4l\��M|��t|��a<��i+��t�b�?�g;i����BY�o ������ȝ���^g����"�{�R�u/��ʜ/�d"t��p�:��#�{Dr?\X�%E��
	5�Q�R0� �N���S1�(Eg��Ǳ�ъk��Z�|N�
_�6�f�3�������8��s��~�]2���^���M�fk��]Xx�>��Ӭ�6 �``���A�u+{����� -N�}��"aNh�J�%`Z4�QcEi��_C�%\�A�Ǳ��.׼z��e�@[�M�x�݇��6qt�L?������N鏂�i��L��R(Y��!�����z۩3(���/�O�/�vw%l���X�<�<�XlxVHYEB     400     160s��^+��uu-̌�
`�pDQ-��VV��"���.,�0\���2�0o&�,���NN�b@E���J��d6;�q���N��D����ўzMmD�&�_R���~���j��F�����'Tg!���O"c(�ڍ���,��%����&����"����-9�D7w4� �ޘ]Wd!��n�#�nE�ˮ���1^ѧ��Gʷ�'������T�Y��N2$9
F��7���������#�V Ⴍ���th>S�ȶ�8LS���:��s��A��c�*�����P^�>1��2�r{j�ϵ�M�용�yl�V�s�5���8p��6��V�Y��l�TlF�XlxVHYEB     400     1408�E�q�; ��[op.�˖�zf��K^?��������0{�[tF�ʲ�^_C�ٛ���oM`p���4qꅔ���]ZO  ������p�2�I�j'���v�@���&Z�Uv�xmA�M"ЖQG�m����	M�R����sZ��7;*ڞ����.�kkU(�m"����-'�������Ӫ�δ�d��H��x�#�fλ[N8�*�Ft�}�n��;��)ic��`LL�c,�$����>��l	Y��B�k���\��3�~��>��<��s�I��ݼ⟏�Ʃ�Ѕ��9�=�����t�bd�F������J��XlxVHYEB     400     160,}���E�,��?�;�=x�Z�1�@z�}[̀�Ͱ�Nk�����InPp(o��l����u������9;��f��\o�W��"S�>�?��-+�x�9s[Q¯gBؖ�j�����\n?�>I4�
�	ۆ�� ���o���he�ӛ1���,ǽݍ�`.)��h·��H�2<E��=����k/Є��	��U����܈Ϫ���C�8ڭ·(d�?�r�4�Ȳ*�(���F��J�vF����;����WV°!��x��엤�%�P	�^�H��#S�g�%\����G�vc���k���\K7+�6|d+���&�-;�;���Ԉ�?4D�2ݰh��n,�XlxVHYEB     400     170{g�2�h�JR�U�7�~c_��=�(sr΀��8�L��G�'~	����'`O�Q��f�7�YA$,�`JY:�!�щ��!��~�	�ի�E�k~?=ݑ����o�V�E�Y��LHv���Zjܴ|U��G[�ҟ\
��(>��R�H�O�Y2r��/�)ws�{�|��w�F��~�2�XV<������O��
a��3�[��ZYw��)p�;�i�4����5[z�9��k�o�c� 	Н�g.t��A���4�$��|&���Xm��҇��$u�bбo�p�'1c-�z�0�>��$J�N/u��d� 4���[�U���=�76���ⵗ�UnK��N�͢�XlxVHYEB     400     160V�{=j���t�D�x�+�����n���|�Ǹ���74�J��2�j��#�x,/�j6k�ҁJ��Z�w�@�v�J�
�^�ִ����\�5����� �t���!3n�A��T��l����5���p|%�l�b	���C��9�\rO#�$dX�����g.3�6��Ce�Y?�rD��TC�vChX���]�h��P�B� x�`�p�/��'l�s
�d�$%"@U~<�`5���x����s��ge%�^�M���Ue���]d��#+��d
t[h��Md'��m>�
�84�i�$UЮ�B�́lQ �|Ø�ۻ��S�b�����TK��	����dWp�(�XlxVHYEB     400     1b0G%i���0n��6�?�P�j�"MP�[�v��]+`�͆�rt�`�:��˦>6@P,ݩ���� sq�MlG�]�]�B�-��::xb��԰�r��'�wZ;2�3R�o�����Z^8D9�H�-��(Oa �� �E�Z��$��#�)�t����q� 2�)�3s=]�Nð���P��b3���]�6"�9���gP5��>=:aW�e�Uo�#ֻ�{Gq�ڶ��G%ڇ� �j
O�,dw�YvgA]���Z�K-���-���?]yve<��hv�'��NO�ӐŗZ�Z0�_�=�C{�Ϲ}�O\
w�v5��S}H"C�o^�}��uT
lRg&���Yd,n<=U]?�����Y�����G�;9�4���5�h3;�0���%��<�Aa@"4h��&:oW�1U�f���¾��~���U%XlxVHYEB     400     110���i�*�O�>K��*'>w���)=��eB�H ���D��-F�(�w!l;	�Rm.Up����>+$ć���(z���r�L���C�횛����硒�x���ýG��ib#�+�ޘ�>[	���
��_A�^��R��b�R�Hp�5+��v�E��C�|e@~� ���_�n6i��d�� 5nK��]iY=�}�װx>�����e�]CT��	���"�'�B �Qn?w�C	�/�ش��yq�^S6�4.%�t\rOg�Р�w��V�?XlxVHYEB     400     180���Tgp��=�$�?�)nu���oL�g��c�M7���$Q��O�R�;�sAn\����]��U��;����B�����Dh/��毪\�h�(I��|M(��G����,�3�v4�-w)�Ve0r��S����F���6_�/1-I��q�j+�����X��ʒV'����e���v���g�o�T�$c�؛&E��*�v+:0�!K��B=L=r�#�j�x��LIX�!�$�)�L���>n&��Tud�ٷ�Aڇ;��hw���E�����,��*7\d!�y1]��:�X1�}�M��M�[����OW�7Y$�fķߪ�7�QYN �4����H)����+�(k��UD��{	
}����O?����UF�EU�XlxVHYEB     400     1800�����L!��b� ����>?d��#�v���m3�jqL���uI"���B8?��67�xQ�E�b-F[� ¹�j�U��Z�T�.J֐[���S��^��V�����=P��`�����wIc� Ej��������_jӦ���2V%�	O^�0,�Nt��F��]m�C\��#��h=��%;�Yz�H�5���X��n�-��A�W6�D635�������uJ�Ñq~�V�乊��͔���1�9?N2�&�3d;��[���x��LrA��	G�6ʈ 4��k�R��5?{�q7�?���6!V����'�S�K���Z��R�����ӈFL1{uu����gV�f��A��=����a	��47��7��XlxVHYEB     400     190�{Nʄ�7�E��:�nA��BRs��8�X��o�nk7��c�jV�OMvٷ}*�g)í�B�`��t1L����� ��
��~}��3.�A��{�,��W&��;q���5����w������B��m�s��l@��E�
Ǚ|�ѵ=�NQIŮ��1�.=��0�m.��Z5�[��f���Xb��֯/jp�~��Z��Z�x	���9 =0;���t�5B�i���"�i���GD���<W�g;r�C�6C"�W��ɉ�X R��Xs�j��(7ݘ+�Ry�Zl�g���=m�=f�jf6�z�+���XmP��~���3������](�m4'�p����u���dxL�y5~t���s���G�Fg+�\��hO7�.i���Ub�X��_�RXlxVHYEB     400     180��hQ:h�ؒ1�G�]�@����>^z�4'ˎ����v?�]"IF1��Y0="i��iqQ�=�u����֧����2fl�[�m��O�Jͷ!�i�ĳ������!r��@��J��R�������A5;`S�7�h�u?Tޙ��f�Mla��M�� 85b|����;���5>K��qb^1�����D�m�H`d�T�NQ=ko	����Vh�p����v�u2B�2�Mz�4@��)�8�M������'��5�e^{T���aSO�z�W<��>K���������H���S&�;�0h�w����/5)��2#W�}��"�o'o�R�MO鏺mJ8RnV�%��Z&X�ǫcύsj�~?M|�O�Z���-�kXlxVHYEB     400     1503��S�d��i�3�ã9y���n�j;%��H���r�'����Q<�M� �0�\�Eb�/ݐ�_PY?߃H�8��êО}�5��/.�6(0��'��Y���x�~2(�Ի5OOUnզ-�c��2�� �L]Ѓ�Z�Z�\��0��o�y�8LnW�T��$����H�DJ�eH�p-�<��X�x/��wC����{��Sr��BTV�B���mhU�5���OB<s})���7����!Nj���R�O6_��n�R)lr�_�q���^�q���}I���̍�h�@}0�,j�O�j6�k_6��@�̮z5��0���'@!+��XlxVHYEB     302     140�8g�{	^��i�q�;Rc&`'f��t5�ZK;0��"�0_e��j���`.�]}5dӞsk�b_}��TA|i��s>�K�l�7Me��U�l���`�8�hJ�7���L��F���<%V�#FO�!�J��PC���E������l�|8~4��cdw*
�ap��}����Z�m��C��E��͠�0��!��C��*.��'4��׷�_�u����9<$�{��3b@�τ�x#�3&�D� ��'ED�$�Yt�p�4��S췎����E��cq濖6�� t�G���٠5��@d�- + 
O��0D�!��O