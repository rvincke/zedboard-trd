XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������8��3�z	V�,�(=[���uu�jϜ�Q��5����>�[��@C:���2��+�f"��J�pE8jC0
�_��ehth�?���@E��y�/)D��^�%D~��m�������)���}�([��<4���O͡ᛲ��A+I'w  bh8mψt��l�Ec�E���������Px�jp�H� :����A˃��iUU;�f}hN��(ti�$V�R��0��0�-;��#��dB�sk�J_Op�,�BHCc�{(U,���!c���]� H���w��v���*�p;���=]^�M���ʮSa*vC�O{��f?��"�W�U���H��s�����^T�?U�K�Ѹ&�7Z�C�XR\!ܓ�fhTa�>'%X���7� ���yfy�OQ�1�M����Gz\ȭ�a�)s�VO��#z&n�`�L�iG9���%!������If�}�`�Z����UV@��lB��*��W�Q�+lWO�Sj-���۸��Eg`q6c���B���Sf��Eͪ{9�X���}�M�eA���.
AT�?�)k@]������Ȼ�߼��5 6�9Ou���ڿT��H8˺�.�q�� \�r�A^9R�2-����s��4nR�Q�o�?����B)r�V�u�5`Q�/�C Q(a+q�k^az�<����_(/�}Q�In�}W�2 �^:��Sc.��g����3�v��s��&t��d��-� #��Aw�z_�y������O�t6į�<u�XlxVHYEB     400     130ȹ��jm����#8=����j�����r*�r+�S|6�b�i��Ψ��5t�i���|WUlKB��b��������(`�F������x{�.��ӯ����0s��C�2yC���*tذ�q8#�5�(�	l�9��:GJ�]b��_P��e[����Ŏyl�n��m��p�/q�v�T��'�Ȟi�eݲ���4���� sp�ˌ���#C�|�����2��u������_b�Aq�[7�?)V�� �ݟk�*#܏xG]Ă�����=������-l}n��^����ƭu�XlxVHYEB     400     100��Ty�iwU�|J(�f?Oh>[��t�-Ϭ��>�Ѐ�b�Ya�qk��s�6�鿞�_���R��h6�u9��{�
x}�I e�c�@!t�����G�5� ^[!���ҜMJ��/bm��I��l�Q��>�PF鍼�b�7�u�*���/wf)�c�������a��%�k�)��ߘ�r� ���enff���W(!��T�E�
�x4	�c��ip����l�!��O���n�bAV-e�ZY�,L�o��#��BXlxVHYEB     400      70�Xd�옼m�A���>BS����<� �Q�_b�qĕ�s-[��t���ޚ|�1�I��0�ýB�1�U%4��o݈۞���%�����e^��;�W���?�Ħ-�XlxVHYEB     400      30��pE� ��o��Y��N�w$t��r��D�0ד�N�X�07���9!�XlxVHYEB     400      c0������In�T<C�+Q�(�S�˻�_�*~�MR���*ݰ5hG�;*}��Co�6u�L�GA�Rc���	�d��N��͙4�XXK0��~/GVʕ;�G���k�P��Z5??��<���;�ܳI+��|?)�Y�˹�$D���U�Q��:����3̪�w�K�Ȩ�ȾV��'���@�O#�0�46����XlxVHYEB     400      a0�-�Nc���@!N��m@�S������G�\Y����Va.��BtD/�T�uL�%��;k����g��Hx�ƣ�~�#��`S���*���]w�eZ����F���lQܦ�e^l�e�z(��3
��6���{�"������<`A��������j�XlxVHYEB     400      a0��(��%}Pc�7X������뮚���bPL���cs@��1E��Ѡook#�^�=��#u���XO!�'l����Z4�!s��w2��f��C]�(ؐ��e�X7��A��)��߈�0���HV4/ 7�NL�BL_�3�I[h�ȽA(-��&XlxVHYEB     400      80��F�����M�`�������x�oh"�*9�kM��Z%��_1���lA�!JC������V�4�Ljw��胴�ր{!=�W;au���x��}^��UHU� ����4|Z>���q��]��XlxVHYEB     400      40&��t;E�;��sw2P�X�����s��i4�����?ſ��s���\h0�;���l�Ә�Bz5XlxVHYEB     400      80^~-8RI(���K���~�Nút��ƶ�A��Di�_ӎ,���ysV�aީa8���\ۍ��p�P��u�|���ѱ�˟	����f���G�cZ�<�Y���Z(V1/�S_W�����[zu�� ��Fk�AXlxVHYEB     400      90i�F���0�|���}����3����Ӿ9K������x4�L��7�ܾ5��]=��ė*ӟ893�;�É}������=D'����
��/29�f�=��q{�6���^G��Rt���R��;˨�LF���F�>�Ջ�n|u2g��<e��XlxVHYEB     400      80�����p��T7��GH\Z�v����D lK$Z�Cx��
C)c��fC����nG��b6z^���lI��!�3=�uf��P�z�u�$&��vA�� �z��  rq\���+^�9�ȶ��xIW]�cοXlxVHYEB     400     170�٤G���ְ���p�e���&)�=�g��xn�Ԡ?�� ��\����`�}��П�ʹ\��/��-i���}68z�"�yKndx��mr�f���a�8�䑎^�)�y	2�0FS���ٗ�Xj��Ň�	%���������6#�+ܳ��-�Pj�%�t�����:^�s������Q`o�F�#I�X:��:$Dp��.�[�Cl���c>%P�+Jց�I���#/�H�.*L��`E��BM��ڏI�#������Lcڴ��m���@������.W��̯%�YYr���}�oo�E�D��@��%p�I��ַ�������Fܙ;���Gu�+��#��V�'��~��؞���
�jXlxVHYEB     400     1a0�.p�O��'�YF�*W 
���Zs31Ahњ$gD	'�?��K�-u�<����1y�ﵺ��D`"F�A�&��h���˄�>*f�wm�uUo-Pf�MvAM�`I���,�գ7d��t�.�����;d�Z���Tr�M�|�s� ���s'�a�Erh����90A�ﻶ�[�G���*c����i�x�g���{&�y��~6�FR��(?f� ����3�G1�T���V�ڼ���V�.|(��3u0m!�-���,G��a�(0������bĴ�*��h�F�e:��ݢv���`��O�ĥ�����W�K����#l��P����l4��ۙ�:��T�ӟ�ۻtW(�OE&3<0�z���c>EQ���+�	���Y\ikaД����5�k�Η\�QC�XlxVHYEB     400     140�N5������N���U}޳��f��P�0�ZH��/����4{��7��K�2x�ϮE;�f*�1�P$���z���@R�>_���fG{�e��/\�|��^Q���b����d@�Ǩ.6j�>�UI����P8{��c�GxI���q>c���3p3	����s��5�6�,O�e��Q��~f�:;z���4v^P���"$1$yb��}jATO7\%|Ju2A���;fq{�4�|N����������{�#K>w!�فGг�ń����ȕ�K�����O�~dH�0��TI`��u8���,��\���XlxVHYEB     400     180gޅ��j?�E Ou�2�S�ѡ3�ޜ]\�`1'$L�u�S��;����M!����v\AB��=VKe G�6��2I������"��]����P�9K�B5@��ohF��䧯�*�CW�������b^���]؈���7�BP20����g\j���ɶ��}C����� {�����z�8�ݔ�_����y}����b�7���?8�e>�Bi�b<�QZ�_��I]e/"�����e�O���1|ՙX�?���p݆+���1 �q\�rTc_$�[a�H@8�����|����V>��K��=7?���R�Mvs�Z���a�ɶ�t��"M	�C�Q�^����A,��x����pH����8�8y>S��XlxVHYEB     400     1b0�H@)F�/$�E<�"�F�t�=���V�J6K�m�K��.J�H��$����3�+�;1�ِP|{&�ofR��W��\ᶒ`!��������&�r3l),��r|�b$��Ý��Up�.=�T{?ER-�d���0�Z'0Y���[��)���N���{P��S�c����^v���iU��:��h<r5t�k����S��_�w�����>|�]Ha7�ĞA���ˣ}l�h��g������� �0�L��u[214@�}�v(O%��s�iJ�B~��H��_��L롋���o���� ���gnyƑ4�؀��7���U�o�gU$1$	�,_W��z�Wz�;�[�`�F�8)���v��[;��7���癈��F��ؽ��/ȲL6u��Viw4����\����o:J��<��{M[�?5�t�ZcjXlxVHYEB     400     170������m�����Mڏ!���^!	��SW� q��]Q�J UU�g��Yk�.3�j�*s_&��W�!N(��s�ϥ�����ɤ���H��>'��l���'s�8'LW��[�L�01�����%�NŹ8��.A��	������'�m�=�A�bh�K�V����0�f_���n����,07��Pq9'��A��xh4�t�!�n�5m�6��F�����1�Mž�=@�젗����Ys1�ҏ�eY���
�h�������ϩs������4��{A�k��ҵ��uY$�\�8���8γ(X5Bz��\��~=Auo�z�LTu/`�~�0�P��?u��:l�,XlxVHYEB     400     130�!.��XVW�����=$��X6�Vr�A	��+��H<���G�^Xo`�0�v���fk�x噧�)H;�T�F�<J��2i�UpF�)��㓂\],��X�B�"��i,�L�Gnn&���~��=@&y���͘�+M���s�8��Հl�|ҩ	PZF4���D����%�L�I
�Y�]�P�����	O?����qS;v����|3����n����.�?]����������ۤt�}�ۡ�E�뭚���m4ŵ�C:���ԭMl���ld��`��5���F�f�XlxVHYEB     400      a0B��DVkC���>ڌ����A��ēt&�~��8��aKy����kޔa�4����ӻ!��
������њ��)b�Dco6*��"��RoD���V0a�kno�0:��a$ƞȀ�P{���\��I�̞��*g���?O�� �bf�b���jbZ{4��[�XlxVHYEB     400     190���46(s�U�<8��Â}P���MR���D»]1����	�-��ǃ����]bs6/�q_q	t�}@�Ӵ�������N1m�ko���F�F���6��'�<r�C���0v/���o,��u\�
c��$o�x��<���j}B)�Y#f���_`��C�F�QI�"��3��4��H7�y� Gs����`�D�(ND(���ϊ��i�W�~{�gXi���Q��t��ܮo��7����r�q�C����F��i��}b8i>��ɬ�9��/�:7�y�~+��hp��Д��c��~��)ZU$.������]�n��[G9��m@�BcJ�����_�V(d�V�p�Xɍ�׈�s��Ʌ" 
�z6eoMzdZB�*�GЗVw�4h��c���Z-EXlxVHYEB     26b     130��6����#}c��6����3"3r�m$���AH̛2� b�[=�<3c�%���4 ��E9I~}zG
3%/#x��w��i���wF!�����?��IO5��Y�N��G����?��#:�j�L����A�ĪT/������]���f�/X��~v���L�YFFT�{�KY�ۣ+\�}y����3��On��`�c"Vk�nPB��cR�.�d󝟝�KDD����I{��:�T�MU.7�ʾ������.l�)H� ���B����ڔ�+�V+�ę�p2T�{lh�c����