XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������2�#���}:���:P�'��>�H��LPU��t�Gr.�� s34�l?�@Z��?�m0���s)�NSJa7Pb�!WLWQ�������+�s���}j^ćN�G,l�m{��L�q��، .><}�q7�b���(��3���e	��I�bXu��R��ֱz6�����^��J��/@���uT���M��Fv1e�Z�$Q!\�+��`~�̧9��`� �^xV���-j�t�xv��}��=���;�̆�g�D0��k����(��헳�Xj|}�rk��sG9}5,���)�,J��}�hl�럑�U��L/ ���g�c�DGZɄ�4vder��^@�����i��
f�����.��&B�D)d�������Ŝ`y:�L��9ʏ�[GLH$�������t]�F1�N��u1z[�#�"�Nyd�T���}=��@��e�u��tEL��	!O���HR=rz������-���n�W&��b�vw�<��.(X�"xgV4���Sif�UU�ü-L{"��?n�,�K�O���N��~�ٟ��ǀ��ASu*4���>h��d�Z��bT.WA�hLn��F�Uqw�[��d��o�� ���H���Ht(��޲�Q̙P@v��G}Ѳ:x��_�/_��f���ݻ[�� ,�EM�f�ڬ�?*S��޸�F����)qzJs{r��$#�.<�Ք��N��ֶ���2η%�U8��H��mOd�[ǜ�l��07	�#XlxVHYEB     400     140�'��=9�ps�|Nsk���턿�"�nY��o�.��P�f�,�@�H�)}���j����b��^_�Y�����2�;�3���EMs^dOSP-鯠/s��:Q��>¾��.�N��9�]tz{��9�f���ɀ�����}�I��{$;o�+X���dI���)��b9��6����&>G��I4mh�ĄWUF���w��u��r����HR!0`��KA.��c��X���]����O��#C���Q;�����,��&\�cp2{?��d��)�y���*z�	��X����L.����'C��@��\�@-Y�XlxVHYEB     400     1a0��|��1�y�등�R�oA<��V�O�����p�	V|�AfN���͞1���1^�ֶr|���ӳ�`ۉ��;@�XF-"d�3]:M=��(q���O�g�Pѹ� �yQ��v=�h�2ymy�P>2���H+A��P���}�0=�VI��P��j���yЮ�����ѡ"�$�y�扻ۂxB��;�QOFѠ�3�o�3w�4��^I�����m�H;.ԡ��h���Ŀ������Ȣ89/ҝ� �}?OE��?�a]}QO�Gٌ��-0
=B����7fUQ~�]``x��������uq� �,ʈʴ������0���ܦ�G��(9��%~CjU�r8�Xԙ%J�$�����wfm��7��''_���ͯ����a �m�G8����ȇۑ�y=��m�I�*Ԣ��XlxVHYEB     400     1d0bi��7����p�}��4�{z��A�!&�`ƌ�9܏t19"f��'W�I:0�΍l���$5�p�j�nk��*���H1t���_�z�a��߳���;��{�&��q�ߞ@���2��P!؜��H�vՇ�5 �gb����R�u(o����P������]�B�A�o�'�kucb��A�6� ��F��Jma�q}�]��Xd� �_|�U��Бa���Ǽ<�6Aϋ|��}��*�5� �*rǶ �����F�t�w���
���4ja�'�'0�S�2������ߤ���{�?x-��ڢ�j��̙��t��KcGl�LQc�OM�A�vm<
)���.��7-©�A_w��߬m!�r�J��V���ų|�w/-z��l\~GH4S
�g��K�e�HJ��#Q`�#囶�k�d� ����-�~6�C�� �I8��U5����t���Bϐ+�L*XlxVHYEB     39b     190�tk9ϲ#�ƾf9�|YP��H�q��0��#"�D	��}�e2�$r�O�-���+rR�\�9�e��� �������6�˕u\��1i��q5�߬��Ӂҷ!��9q��D޺�r�@������hh}.I����q"�e�-Ț#*:��e�|e#��L��}a?��nF숆r
I��}c�+�䵌�;x·��x��g�����I�i��߇JYL��kZ�Kr���YU@�&�Hظ�ad���X�#�ȶm�j��K�%�\\��k�&�D��EY�X�-Ȥ�rJ2:����@n7_L@u��- ��Fvx��J�E���J�V(A�IK�<�qE�.\c:4������6�0c��f����29�c�ُe�븾�}�~r��σA��_}Br"ӮL�/