XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ߒV�:�d*گf:В�v�F�wP����� j��:�*89f��E�$u���d�#�ΈZ���v�˪�����@w�~�]���#��ظ�����U!G?�-zJs]���M��6_�[��'3�xQ�W�)L����F�C6M^�r�]��
�6酾�}��9���`;�y���1�h�ʰ��ю��ʍ	(�I ��?e=�ñ;r��^�BIY�ȱ�@g��.3��4��v�q��{b:���ެ-���,�=��f|5`]bg�(����#¿�0�&(��}�X�noP���Vˊ.��Hh#�""�1{��,�;(XѓѴf�_�1�$f�皏�0:7FsfVj�r����1� ����Ј��p�J*]Slzl`��Z�m�K������v�4��<�k�������hک��
Np70L�@/
��\k�:� ����6�.���w�Vz'`CP���� =w�կX�`����fo�{N5
�q]�h���%ؒ�9p�n�������M��1k�3#~R^��]�0�����w6�ҭJ�&I�p%'W���<��]+!J�Jz�K��ߞ�YS��lgڑ�liݤ�
�Mp;�%ȝ �E�}x��bN�%!���N�ȴ��|N�d���L���s+�é��s�"��?8D.��m)�6��ө�}�ca��;v�d.�M�h�
%v�Dա� ���`�����:�d�7&����'ؗ���W�}n;<.j���,�i��;�nSXlxVHYEB     400     130V9Q��w�h�������4�榥>.��cr��{�u���2	YC=�����K��CL$��8���n*�`Ӕ#B���4�&6R��F�1�������{��q�L0^f�(��0�Hdk	)�"r�Q� �گF>�84�;���E�mˠ�I�
�D��0C~~��XLU-	��E�W��A^ �RS3��OM���'����I�M8���Fq��5�(�N$OCrK�>Դ[�G-�%J�KB��Ys#��6ʀr�Sn��������;�����/
x����7Zm�:�qU�k�ӫ1�J0�hXlxVHYEB     400     120�3�j�(�(�4�h@�=3����_p�(x���bXʀ��w�,�?P�����m��j����l�M��d�O�{q����]�K�O�}�'��`I���)����ȕiv�`*�l���c�x54O�+¹�SX7���������3ҩ9��{C� �`���ۭO��oW|�q����j�90��^��tf�E��Q�M�ģ�U2%h'�!�mi��[��}ᷦDA�?X����������� &�j:&
�������2���l���!}G���@��|= �XlxVHYEB     400     180g_`#����������l�ih�x��b����>
�H@��O-�dП�����_Qg�lŉ� '��Q�*p�V�&���J���Y%f�͒���럮��`����j&9gf�zyv}:�U�Dɨ���А�z�bY�*>�{��np��Aw�W댕�&y|��s��m�&���M|s���$�q!�����#�-���2:����˱C�_����m��v�aA$�LV|,�Kn�����@��u�ƑD3J���=
�1]1��T#��k�D?�mا�?��e���(����"����!�G��o�ʒ�,������� �t]�! �02@�����Ĩ<ds ������
�8|M���eMM�5� �'��w�Y�XlxVHYEB     400     110Z�F�7э�3��~�M��'3]�u9(UZ�W����rj�d�v�6X`_F������?D�ze{ٚ�A�j�ڇӯ�I ��)=v
Lv�D���_i���l�aL@b4}Y)e08��2�L���{{fa˛�@� <�K�5��z>^�B
+�Rv>}�Ubw[�}9�������XH�w\������ 5�a�&U��7�S7Gis�@������\�/t|#ItL�j�E�M�I�pHcD�ؠ�Y��z�݅�[��SZ��|9XlxVHYEB     400     110���f�g�����Z��eƷC��ezL`�3o!-u����'���ҳ�`%��EV��tח��m����}p�3OJ"[g��fx(�r� Z��̈́I�H>��7�-�o�ߚ����Ԁ�&�����S$˅��>_H�ܸ<��uP�8b�<l�?m����"�e�$�п^��(��@�٫h`���L��䵂D.J�<D�]�V<j���=�A�������CUH�(���<�V��R=�7�;!�\{Ӄ$��#t��ܺ�L��%zd8b[FXlxVHYEB     2b0      e0w�o9M?2$�{f�������@��@��zy��e�u,��!�٠��F[�8���|����Ĳ�o��^���"�q��M��F9W�34V���� }~#���孞�|�}�l2��9V����V.h�+��HU���᷍�����n�B�၃��_`ӷơ�������eB��G��<r��[��tT��5ʌ��	�J�ܰ�QPv�|������.l�,V�:�y,