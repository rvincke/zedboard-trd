XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6"1L(��ޠ�1�Tw�YI�m����2�w�J{ �Z��ӚV�9o7��}�[as��Q��hG�K�g���8��2�w�O<�R�L�_kg$�	��nt��
(��E�F��<�Wͯ�w��:ƞi����������
�Az#v�ɡ�������hi�=�F���1)�@_t�Ĝ�@��0.39��ʍ����	�v0>��GΊ��De���[��T��6�R=��Ao������zC�N����o2$�}m�j+U�^�³�\�I�v'�����Vt:-�?�Xr 8Nb��V7{�fr}	4Ͻ"�y���lPzw�0�����@���w�	AO�o4�?5xO�u�|�3?b�&���Nu6!��8TA�OѴq���2k���݀Ŧ�/��M!�PcY�܆̀v'��l�H�_<��eEх��=}�5�9Ý�'�*���k���C#H�0Mw �k[P�X�7�X400rj�g�w,�����OX���Ң��nYiK���W��p�G�<(�(�1�!�F�]$0{Z��F�t��	ʭTy�?wA� ���q�eA�����U�%]�#�gY�zG�M� ;��Yݹ�4�^׾�#,,p-�I#����� .�\�]H�X�b8c����ђ��T�\�4ߵ�=�L�� X�Ki>���ZX��xKY����`��R�o��8�<|7�4p�S���=���Q�J8��(�"����gUl���M`݋��<���|�!���M���-0?�_ݬ9Юn��ۈXlxVHYEB     400     130ю�֦6^7L���
9%	��9f��X�EI30�J���hS��9�"� ���U�lB!s�8B�˔(T'�\��m�%�� �×E" � mP�q��@n����W���h�U� -��H��Ď�1��`�q���?
�O���(5>�J*ˍ?���Ⱥd?����;��6$�A�"�U1��!E�c�ǿ��w��e;�=����%���dK)%���e	'q�����`��`�\Pej$��|Ʋ˦nY�?��_Ko~�3�,�:u���/�\/��MD���]�5y�����iM�N�XlxVHYEB     400     1c0܌�;��XQ{����AÎ����ym^b�h@��6���>j�9-D��a�8���ݯ����˃wYN`l����{�x�BU�}*��D�(��+L��(Ǚm-C8�KӸ2߫������
�b�f�2Ue���1tș��֏��JD>�W�&���C~��D�z��-N!��ίB$^��j�A�,DHR����|ָP(�X7iヶ$�a��l�a9�戥*)�m��:j� .GM �����Lp﷿�Ku
��tU�5'C��}���X(���t�������~�]8c�5P�:n�?���<�wu��" �s��,g��&|� �V��"�*1�W�����h����w�1�����I<C45�x{�������;:^��6�Dp��h��Q���q)�gPo���}��/X�+��P���}&z��fj��{�F�XlxVHYEB     3f7     1e0�)��BS���@Bް6�5�	�PjU@Oxɹ����kS���`�.!�*� ��^���ur6��F�7��xsG�zƟ�S�N�AmF32��Փ�=���v�)������Fɪ�$A�F��e�-�\�3�㙆�J�.qtP���W��J�H	6���y ��(j����k
���xj�eHߜ��;���a	k�h�9�3�2*GMlɫf��6��O��gS?X$ɠ�z¯�]��p�߽K�;}�x�֙��x��$
�4��1�����~�,�1��P�4���x�3���}˶�����kM����a(����S��/>�*�G��=i��n6����	��zg2��#�/{�3q5�ʮ�qȀ�%�4�{����nRٗ���e���dLb��ΥX��oJhӹ�7��crhn�`t��,�P�-���R��^�wX�k�}�sf�Ȫ��Gwyx&���8���hj���{����=>�