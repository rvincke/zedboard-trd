XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�~'���o[�C2���
0y�;�Y>�&��\�%{�����K�1��0m�gE��p�z�t�!�_��-��]п1R��]F�8�o����:��h{ny=��1��Ó�O�3��:^���>y�	�B�&�W�#��	bU)4�)��2���{�{����`�@C�����#�.*t�E<��k�g-�5���Q��q|��Z�j`w�}�HJ�v��g7����c>|E��w7�E�gݨ�!5��A��0���i|�zO����Ʒ��'�L9�a�;Y��3�<�:[p	�e�D���iח�Z����k�Q'�.f�110�j�7�|[E�b���I�U�?!`�N� e�2���QW=
��V�u�HE����7'��#��q����:ǆ��+��`saٜe�T�����w:���V�K�:n�6ҍ���E��A=d�|��/=5�G����������9'��كi��Ly��\�w^��ŵ���{�&�i��@޺O�'3�����V:"����:W�YyӁ̯Ćv&��?���C��~	�����f9������`5Mg?��~�7���y�.wvA�� �D�����S�/��������0r.�|��,�ڒ�S�����_B��ʖ���=�A�8V�`�Ύ����0~��,k;�1����"g�i��L�LfR��}`���8mW�F��φ)���*Uop2	���0 ���[M�{SLv��3��f?y���GE�D�2M��Z�0��EXlxVHYEB     400     130�j�ά?�S�&�kks�0A�m��e��5���{B�Ղ�֊�q�S ���iH6��HA	��xW��hA6WN�y6��=ʀ׮�i4�����#�W0��>&I3�lw���
�T<Z��G�h����"M7����Fay�+�N�Ms��E!��WldN�g����X��]�7�1�=�C������o���Dg�z�<h��x��k�� -e%P�BTg���H` ������X}6ܯ�C	��@>qIg�㶣�Q�g8
��]���С�Y��o7{���SZTQ��?�۽�"j�XlxVHYEB     400     150��d�_�J�RA��-tL��&",��kU��cQ(�cc��u���[����ulD��sc*���H��}k�P?�'L��37�\@7���7��f@#c�9e���k?S��ͭ��X��HBqx�e��1��b.��x�Ox�r&�++Ц�.�]�?�ҾF���	>��# ��+����N�u��8��^�%!�߿��AKT�9�]�`ilX3��� ��Q�]�=?S_�Iz�!]�˟P�&4U�����5�}]�����݌эo���"Gn r�?r�׹�a��ɚ�c�i6�4���?�q.��Գ�'�Y��|�F'��ۂ���XlxVHYEB     400     110�P�+sd�'��*r�懁Gi"#�,�@Y�a��b�bv=�o�交�a� q�F�>u�����ܽ���>5��&陧,���?�����(i�}9�kO�i'�yv��~���|���7#P��蝾َa�����X,��t�Y5��:V9�V3#F+�4Fp�-C�熭��z�*�Y���%m�mY��t��:9�^��9e�4j(-��I_�����u��6'�2������'G�)n}� �I��0��R��� njjI���t���OjiJI�XXlxVHYEB     400     1b0��)�\&�mG-��w
�T��9s�@���#���4a�`�vh>|�cA��L+8p&�1Z_!k��e����z�9.���6��5t�%��-��"�I�����ex��Iz���r6�ŤBMn�7}&Lz��c�{�n��TK���_r�ɓAH�#�ק>"f-��I�'������ �y"�rE��~9p�8R�0z�CW���>�L|��O�K�1P�L|1jq �n���#���p�G�3���!���h%#	vȌ���P������g} b�'Ν7���������p�:Y�p��ج�],�Kٸ�W�p�� #�A���cY8\.x������N4����4��G^��%��+�}�2�oyn�mwM�L�;'��
�*bJ£�Rˮ��(���L���/G��<��T�?����{XlxVHYEB     400     190�Ş�G�B/cd�zX��:4��Ns:wm� ?�36_��wsD�PgDs�,W�wo	��6*�w�v�3���W����7���{��:gn�Q� ��BX�czt��[���G"$���.eJ<�&<��90{Ҹ���&�VӮ*g+�B�u�!���������-?���c�hG8�`O��c�{�|��.���pP5C��V�Ǔ������-�Z�����	v �kW[5I�;I[��}��{V��C-\r)��~�C��|doW�o�j����c�0�	��0f�`�e(I+�e��2��ܧK��o��}��iA_jR�������[����7j
��)�*���.�M�Os������e0������#�Iκ�.���Bws�� �m�	���XlxVHYEB     400     150He�������Kr����m�h�EeP�~s�"_�E�Ě-d�r�%d�><c=�=ᝇ�C�{�C4vQ��An��즹8VX��^jY��c��������jf�,��^[������\��b_Z�D���+K���0(`:B��26羐��i����=)<���7�	�={C��nK<ޛ&à��ge��f���yom"	:͖�61��3%ԪUn���seGvdNp�+gV2�v�E�Q�U���5.�	��CZ�!��v����:6Y>��\����:�`�ϡ�:���}��gS�38y��ؕ~���Ʌ4�&V�v�	Rt^��XlxVHYEB     400     160�i��n=1��#���I�>ئA?S�*�"V��f���W���r�s�̺E�3�.�S��\��>�%��K{ǘ��ni���G<?-�m(ؖ���UWJ٤4��U��5[!���=mC �;��\q�v ٿ kR����\�?��c���՜6�8��b���1�� �*��B�,j��8�6�w���pIY�
��.;�*����Uw���7�;S��e�����ګmSxY�1U�D/�%�] o�$�[r"�J߮�S)
���Q�B��f�M�	�T��hk:��0�}��Y�Ď��r�#L�q��l��By�_3�Ձ�}�����f����ͅ���Ꮪ@�>[~;���y�XlxVHYEB      7a      60�� ���Z�:�O�W~�aʡ,���iؕbNU;]����CIȂ`F�L˳p�&�h9]̹�P"�N�}�G��b[�7G�2rj63<܆�D�*�Ҧ�