XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����J�,N"~O�+-��e&��\7t*	�C�k^�ۄN=x�>�c&�#,m����>�s�7�����#�Q���P�A�/z�Ɇ�w�P�?5b&�f̬9��.}F~��jY/$K)�p ��=.d�Q0�����+�W_fZͨU�� �״�#�� l��5f~����2'~R�"ile����(�JR[��7���7b6ZU.&qn�6��XYߜ��g�R�I���os��(�g}�P�llKX��Ff����Ԗ��5y11�*�2�@o��d
6�/:�����N�j�R��б>�)��ݖ\�D���v�=�@���m������7��6?k�63�I'-�7���@9��K����\�.�W��
�4�s�Kt�ӻ�\Y�N{nI��پ�H��<hL	����5cE7m(�!D��>D��F�V!�.�3����N��4W7��� ���e�Z�8Ɂ��?ZR�ZA����L��GW������ 3�쀒Nク�
���p5�	iz8`h!f�Kp∼R
�GK�o�:���$P9n+ᵢRn��Μ���Z�`�j�Mׄ������̝�c9GEu��dq�r���AD	�ʤLߓ�a�͖�ОY�l]۸��5k���:��o���ʹ���lL��g��b��j����eX����
M�����g�@�PV���/��rՈ��xg����EQ��R�vg��ݏ?����� v�B��הJ(�Eb��B���tׯHU��	(XlxVHYEB     400     130n=� q-֌T_��m�~d�
lT�%�߮t�y�@R�&�W�<sVp��:K���Y��>�/��vn���IDQ���g�M��Y��"�/:Ş�|qOk��%���Zpwgx^53�DIW1���K�xW��������^5�Y�p럭�tg]�4��1�T���v����G�M{�p���8�$������qq�Pޚvǳ
�� N�!r��k�P�g�S�=Cq�wl�ڷ��W��i6/����nZ��~��w��]�g�r��-�Y�i���1Fo��s��ZdY�RXBN̚��� �'NLXlxVHYEB     400     130V���,��@�wL��#�^�J�{�°������:{!AډB�K�&��1 ߌF�6Qz��ت�7q��x��2�?�U&��7� �8��u��0v��O5�Q+f�*)���)�^�X㰅{ޖ��5�:EOB+�񧳆���������(N� A�GLHY�L�=yM�}G�?s�`~*�uI���e>ЛF��s�P@�Y���\y�Q}L?Yo���n���R���E��ZO�=0Nv�gȅ�x�4	���Y;Xg\�K-�$�~���'��,{8��V��F ߜ�|Z�$ǒ���D�vej��<XlxVHYEB     400      c0� }��U�L&��?������$��j���W�'��9<R�S������P2�K��m��5U�I�2�8"��)����j�����);z���;�ݢ���W��Ŵ7vN��E��FB�$ID���@���͗q���N��D��K�	��:eBa��>�M���v���>T�]��#XlxVHYEB     400     160�$���dY�u��2�4��jLW��5��H�:�3Q.�}$#Ҕ.y�� ��364�{D�����I\g��3�����v��N�>��*P�MS�v�@�`��PphWr��������I��~�*u�R;���t^͕ח�^��f0Њ�Z~T�%��7���y,�dy��%_%c�ď�-�ϛ��6���� �>��'Iyc�.g�������0W1xE����v�V3��$�TW&Ҹ��
ڜ�ze	X�t��;�B��/���
��I6����rȷ%f���Ʒ3�Iaf��gP!@0���9�.J"u�c[���%P��7a)ޑ����.[G��A�Bc��Z~��>XlxVHYEB     400      e0t[CV�X'��H�?�&rl����7�q�����i5r�ֈb�w��~��9�>�����A|�0��2�����8����ԧ��H��m���b����	�����(޽Y�g-߸x�F`~1�v�"^j��l�O�l�r���sOfR@�Ϝ�h�N=:w��9uouw���^牾5p/���X!�
�HR \������oFK����6X��߄���S�XlxVHYEB     400     160[��*���u���En#[��j�&b�x�d�r�c�[�ga�_(�z+A����q��hV��<�K8�V�+�(�.z�FW��8(b��\V����H"�bg�Y�T���b,���gS�����(1u1�%�\��D���5����N����,~�^�p�.'���H~���x��;b������^��(|�m`�~��ڐ)���՗��ə�z���i)����30��o�i �<�隡�v�H�(�d��8kbl�fԄ�D����n R���xa�6��:�je]
� ����x��U4'�M�B�n���t��8P���M�b�ؾ��z��G�ۙ�]�����XlxVHYEB     400     150֦M�7ָ�-���su��ܜ�گt,�"��US�=�h�Q��YH��2��DFb��i����P�1󐀖3�U����~>>SyKTR�.tJRWR<!X�{D�G�4��I#��#^J�vyQ�f���R^l���$xӿH�����d~���`�E�����I�ǯ�@אŊ���zR�,�t�O��Lf����h3@�a>�Q��S��R�����Ʀ��}�*,=��!�����i�h��$�B1�j/�;/�}���������brj�ί�M~�PJ�{V��뒱�iz���X�z�=�Ԝ *�\�qc�P�$��%��Z�R�_��XlxVHYEB     400     100j)4A!Ic�bs�(������O >�ʕ�3�žc�pG+��3#>���N�Ĉţ�C� ���Ӂ�}�v~�D��s��S���nfb^�Us�6��A89:�)��:O����B!n5("�T�i���<_����S
7�@G���2	'a�	��J�t`���γZʀ�����Au��k�����[d�p=e=��<1����ퟺ��D;9S�ՐU��$C���"Uڡ���8P�� W0��XlxVHYEB     400     120{����WH�G��7�!��*�+�!�������ήG���:=$0�l3V��{��5H}�x_.�j�m�C��nL	G�M',E��D9]�b�p���Ph����z��짊φ�΢�� ���#J$領��q�����w@�C���:�͜�2���cԀ	S�xz���X*'F�/IW�I#\�ک7�}գ�mi}ܩ��# #�@����G�7m��8W9'�p�As�ۢ��nP�
Wy݅a����\�r��1L� �`g/�~�r��|�Mh�XlxVHYEB     400     150��Z���9��7\iR3��0��DR"^�g�!��pt�mLݞy=!�ם�Zf�~"����<���s����P�̢�H��� ����M����VcZ�/�K{Nv5�h/�����A�% �� x0�:� 	N#�r��]K��m��d����^���(�C�V���f^��+��bo�ϓw��/[��䳟�v�`^
���4,DZ��I5to?���Y�S�_~�cOs��M.��$�;'s�B�H��<lt�ȱGÎDI���>����2�eY�������i��DႤw�:Ϙ�U��z3pd����W�5v�{�Q=<�^xX��z�V�cPG7l�XlxVHYEB     400     100�vp[@�R��$�7Y��� �6��s5�xy��aN?�������)�����M�o���:�]��]���Q�n�^IL���({���,i�x�˅nϰ��Rk��l����� n���)�"��&���Z���_"8X�6�b�W��8X$wV�	��РA��%�,�_�a���{�K��{�(��T���Y�Hx�.6�"h�y��Mֈ/T#;M<��u�Ӄ2-¿�w�������n&������k2?Ș(t����������XlxVHYEB     400      f0���d��Fe�sm�̠�zF���=��Y�#��t�p�]u2����{��c�4c�޲ ����a�qBj��Z�>,�O�!Q�0�]xR�;�$�����T���K̹����gHҎ�&m1��oٍ�I�����b@����u����g���V*�٘�z�*�zQ�FO�A+W�5���;�;��{��!<uH�d�l����n	r�h)�Y�!���F&k8WM���h�"<�XlxVHYEB     400     100ES�c��m\4�{�\�����uH�
���������_7�����g>��jf�ftd˟����4�O����A{4K���}:���B���X0P�!��{����:ǚ* kԢL��=0�#p�r?$�/��7O���!���W[�T��6�v��3�{�� �W�l�'"�G�ۭx�����q[9���9����Y�i����7��j��֓1���q��Qxx�Jϒ<�S1O�����f7ZH$=I�������b���~XlxVHYEB     400     130��;����*� OG�yiv�I���~���a4�]ۿJ�8�:@_��A�E� MM�+�j$�VP�XUpT��c�i�l	�{d�������]����\�B=I�ϔr��@�RR�'�yH^��8i7�	�_�qW�k�%�6jr}/H���wQ������"��o\��A��ʁ�$A�َ�V~�K��ZP/HTGgL+@��m܃?� b@ˏvJTI��}�8��:��d���	�:X��'���o��"�C��ܱUp�UC�\V��I���Vg��� pB|��}Q�����a��~�83kEΝXlxVHYEB     400     140ܯ�ɗ��U�c��E�X���5�SF}4ү��-��!q۔�>�"��k���|ȑ7GA�ř��mx>}�',�2����s��K�u+ޭ��5z�ׇ���Yʀ�F(5�ݗ�b�8f�&"ûɥ&��7���j������4)*&��}r�爹��4p��O��B�ż�,��<?V?���Rz���q����	��$)��>�_%��Y�����"	�*o���q���o6�{�e
s:�(�=xЩ9��?&-�=��a�3 �'i��1��t��F_��jD�P�˖D��*GaA�X�B�7���< �EĠmi��XlxVHYEB     400     110�~�9G�!�
2?v��\\2=q�R�#����ɳ�f�U�����B�t·3{_�<*�]�Ю�ʤ@�-����N��F@�ܚ,⏥-�;2���jEt"���9F�a#K��]��hs	��l�8�9�7�E�_���u	k����@ZL0��\��>
 /���������-Q����E�򊪽l��N��[�̿�΍��b���ѐ8�-�d��1��k@}��*s�v�0��R��<�-z]�.� MP���)$���G�XlxVHYEB     400     100u�6�����
�"���@�)5�E�ƮeN���<��45P�$q��W�G(�J�3;]R��)O�E'붶f:�;���pV�}�z�%�'�=voȺ���D�,�Dk�����Y�vy��� mf��eƎJ�O�MF�f���r�������86�ϑ�+�u�+�Lƨ�`��`d#�ܚ�X&4v���
�M� ��-�C�����7"H�2-���0n���-v�x�� ��M�<��y������(ߕ1XlxVHYEB     400     100HvK`��"i�v�4�����ۆ��Bk�86$��ۚo�-�.4��"rw��V|(ۼ۰Z� �w����x_��T�J��2YEdO͑�F�Z0X�Μz4���gn���Q��U	�����7p�Kdi��l�^��&�X� 9K�Pi�EKȤ�`P�.�/Vc�ؔ�.Ծ�?�4�Е7ϙ�1��=��;JW�@�~y�D_c�y�@X�<ه���DY|:M�����xˊ��>�1-�޽N��[�Y�XlxVHYEB     400     110��b?��+��ǻ�ʭ�|���͛��6���De8����8�$�F9����b����ux���� /=��ӧ�Ñ'VhK���,���'����Yʲd�kG��k�IP��%�O���Z�My�������>q}N���~1��K���B���%1�H֜���f����F_29)Wh�#4#�.c����W�,�K������݄���)2ɋ0�	 3:����A�Kp�	A�D�,�e���		�����xR�'������Z��@�XlxVHYEB     400     140w���6�8��
��1�-�z��39�SEq��T�������Ev�U�+lJ_��3����>N'n�;�r'a 8P���Ɲ�M9$��G�,�g��ה�5�f�aѣ	�������L��§r�-��+�6+�p�H��p;��;�H�L����-`�fDv��8�22��kQ:�mD��m<l�JV����?٢|sX���ě�Lg�#=?�ףi]���)n��[��Y}�t���X��?�j�v�]�k�@iI����K�9�5z��<�D����Rs�24�B���q����̐1{/��7?�/f��$Q���20XlxVHYEB     400     190��fC�g=7�}�Nl�֊��!��	[%f���n%k� �p�� �|	^EG�v]&���(�����5�x�x�r޳I��S�.\�4�&8��~���2u�����,U��Jd�y�$NԬ�ɼ���?�yC9������l��d�w��/��+�eC:�\�.�lSpVG 4Ba2��|=;g9��q	�V����%���]xU����[m��R~ܶ�>&�ق�iʟ�(fd��eV3
���~�>�:�*�)-4{O�G���%�m���=#��i�����f�.���R�}R�rڬ�2�;~|f|��_G�[`|�uai ��Ş��Z.��q��X�|M��	�����uz��ֽ��4��9·jd�_���Vm�ˑT�~��Z�F��5�XlxVHYEB     400     160�"��Y������C��F&m�m��	��-]ض�-��u�dU�0��Xs?X�
�ma�=Z+_��S��=��
�Y��s���u�#�Nc��c0}v�Y$㵨s�����bJ/���v�җ�űG���E���`�I	�"��2�;H��t�Ns�i4�]#E'��Ѭ�x��܈{Z��g�!am� N�L�����QF-����+��uJ7ﺏ��Rk+��M�i��*\�E�
f����MPb�z�׍�:V�E�T~wOF��;ʉP�h��ǑJY���WU�ٟ��_x�#�'�},��M��ԧ�qg�qJ�%3k�����6L{(����by#S�����XlxVHYEB      91      70`�d����>[�"�!�@�#^_����Ո�S���J!���-�Ku�Z�}�0��/[�@�I�`k��7����to�pOm? �,r���ix�1k�&V���,���{�#g�d��